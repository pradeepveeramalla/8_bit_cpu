
module and_gate (
    input wire a,  
    input wire b,   
    output wire y   
);
    // AND operation
    assign y = a & b;
endmodule
